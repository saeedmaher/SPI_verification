package shared_pkg;

    bit write_address_done;
    bit write_data_done;
    bit read_address_done;
    bit read_data_done;

endpackage