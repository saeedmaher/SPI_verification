package shared_pkg;

    bit[5:0] count;
    int limit;
    logic [10:0] keep_arr;
    bit is_read;
    bit have_address_to_read;

endpackage